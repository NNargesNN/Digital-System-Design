library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

use work.Convolution_pkg.ALL;

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.std_logic_arith.all;

entity convolutionTB is generic (i_width  :integer  := 30;
	     i_height :integer  := 20;
             k_width  :integer  := 3;
             k_height :integer  := 3);
END convolutionTB;

architecture tb of convolutionTB is
	component convolution IS
	generic (i_width  :integer  := 30;
	     i_height :integer  := 20;
             k_width  :integer  := 3;
             k_height :integer  := 3);
	   port (
		clock:in std_logic;
		img  : in vec2 (0 to i_height-1 , 0 to i_width-1);
		krnl : in vec2 (0 to 2 , 0 to 2 );
		new_img:out vec2 (0 to i_height-1 , 0 to i_width-1)
	  
		);
end component;


signal clock_tb : std_logic := '0';
signal  img_tb : vec2 ( 0 to i_height-1 , 0 to i_width-1);
signal krnl_tb : vec2 ( 0 to k_width-1 , 0 to k_height-1);
signal  new_img_tb : vec2 ( 0 to i_height-1 , 0 to i_width-1);

begin
	cut : convolution GENERIC MAP  (i_width   => 30 ,
	     i_height   => 20 ,
             k_width    => 3 ,
             k_height   => 3) PORT MAP (clock_tb,img_tb,krnl_tb,new_img_tb);
	clock_tb <= NOT clock_tb AFTER 10 ns;
krnl_tb <= (
          (0,1,0),
          (1,-4,1),
          (0,1,0));

 img_tb <= ((255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255),
(255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255),
(255,255,255,255,255,255,183,32,0,0,0,32,159,255,183,32,0,0,0,32,159,255,255,255,255,255,255,255,255,255			    ),
(255,255,255,255,255,183,16,0,0,0,0,0,8,120,16,0,0,0,0,0,8,255,255,255,255,255,255,255,255,255							),
(255,255,255,255,255,24,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,255,255,255,255,255,255,255,255,255								),
(255,255,255,255,255,0,0,0,104,255,135,0,0,0,0,0,104,255,0,0,0,255,255,255,255,255,255,255,255,255						),
(255,255,255,255,255,0,0,0,255,255,255,8,0,0,0,104,255,255,0,0,0,255,255,255,255,255,255,255,255,255					),		
(255,255,255,255,255,0,0,0,159,255,255,135,0,0,104,255,255,183,0,0,0,255,255,255,255,255,255,255,255,255				),		
(255,255,255,255,255,8,0,0,8,255,255,255,255,255,255,255,255,24,0,0,0,255,255,255,255,255,255,255,255,255				),		
(255,255,255,255,255,135,0,0,0,32,159,255,255,255,255,255,183,0,0,0,104,255,255,255,255,255,255,255,255,255				),		
(255,255,255,255,255,255,8,0,0,0,8,159,255,255,255,183,16,0,0,0,255,255,255,255,255,255,255,255,255,255					),		
(255,255,255,255,255,255,135,0,0,0,0,8,159,255,183,16,0,0,0,104,255,255,255,255,255,255,255,255,255,255					),		
(255,255,255,255,255,255,255,255,135,0,0,0,8,64,16,0,0,0,104,255,255,255,255,255,255,255,255,255,255,255				),		
(255,255,255,255,255,255,255,255,255,135,0,0,0,0,0,0,0,104,255,255,255,255,255,255,255,255,255,255,255,255				),		
(255,255,255,255,255,255,255,255,255,255,135,0,0,0,0,0,104,255,255,255,255,255,255,255,255,255,255,255,255,255			),		
(255,255,255,255,255,255,255,255,255,255,255,247,88,0,0,104,255,255,255,255,255,255,255,255,255,255,255,255,255,255		),	
(255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255),		
(255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255),	
(255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255),	
(255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255));	

END tb;